.title KiCad schematic
U1 a NC_01 NC_02 NC_03 NC_04 NC_05 NC_06 NC_07 NC_08 NC_09 NC_10 NC_11 NC_12 NC_13 NC_14 NC_15 NC_16 NC_17 NC_18 c NC_19 NC_20 NC_21 NC_22 NC_23 NC_24 NC_25 NC_26 NC_27 NC_28 NC_29 b NC_30 Net-_U1-Pad34_ NC_31 NC_32 NC_33 NC_34 ESP32-DEVKITC-32D
U2 c b a DS18B20
R1 a b R
J0 a b c Conn_01x03
.end
